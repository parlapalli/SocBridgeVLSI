#welcome to socbridge
