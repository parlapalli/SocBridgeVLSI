module test;
  initial
	$display("Welcome to Git Repo");

enmodule 
