module test;
  initial
	$display("Welcome to SocBridge Semiconductors Pvt Ltd");

enmodule 
